package Ram_shared_pkg;

    parameter WRITE_ADDR = 2'b00;
    parameter WRITE_DATA = 2'b01;
    parameter READ_ADDR = 2'b10;
    parameter READ_DATA = 2'b11;

endpackage : Ram_shared_pkg