package SPI_slave_env_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import SPI_slave_agent_pkg::*;
    import SPI_slave_scoreboard_pkg::*;
    import SPI_slave_coverage_pkg::*;

    class SPI_slave_env extends uvm_env;
        `uvm_component_utils(SPI_slave_env)

        SPI_slave_agent agent;
        SPI_slave_scoreboard scoreboard;
        SPI_slave_coverage coverage;

        function new(string name = "SPI_slave_env", uvm_component parent = null);
            super.new(name, parent);
        endfunction : new

        virtual function void build_phase(uvm_phase phase);
            super.build_phase(phase);

            agent       = SPI_slave_agent::type_id::create("agent", this);
            scoreboard  = SPI_slave_scoreboard::type_id::create("scoreboard", this);
            coverage    = SPI_slave_coverage::type_id::create("coverage", this);
        endfunction : build_phase

        virtual function void connect_phase(uvm_phase phase);
            super.connect_phase(phase);
            agent.agent_ap.connect(scoreboard.sb_export);
            agent.agent_ap.connect(coverage.cov_export);
        endfunction : connect_phase
    endclass: SPI_slave_env
endpackage